module cpu();
endmodule
