module mux_4way16bit_chip_tb;
	reg [15:0] a;
	reg [15:0] b;
	reg [15:0] c;
	reg [15:0] d;
	reg [1:0] s;
	wire [15:0] out;

	mux_4way16bit_chip mux4way(out, a, b, c, d, s);

	initial begin
		$monitor("a: %b, b: %b, c: %b, d: %b, s: %b, out: %b", a, b, c, d, s, out);
		a = 16'b1000000000000001; b = 16'b0100000000000010; c = 16'b000001111100000; d = 16'b0000000011111111 ; s = 2'b00; #10
		// TEST case 1
		a = 16'b1000000000000001; b = 16'b0100000000000010; c = 16'b000001111100000; d = 16'b0000000011111111 ; s = 2'b00; #10
		// TEST case 2
		a = 16'b1000000000000001; b = 16'b0100000000000010; c = 16'b000001111100000; d = 16'b0000000011111111 ; s = 2'b01; #10
		// TEST case 3
		a = 16'b1000000000000001; b = 16'b0100000000000010; c = 16'b000001111100000; d = 16'b0000000011111111 ; s = 2'b10; #10
		// TEST case 4
		a = 16'b1000000000000001; b = 16'b0100000000000010; c = 16'b000001111100000; d = 16'b0000000011111111 ; s = 2'b11; #10
		$finish;
	end
endmodule
