module mux_8way16bit_chip_tb;
	reg [15:0]a;
	reg [15:0]b;
	reg [15:0]c;
	reg [15:0]d;
	reg [15:0]e;
	reg [15:0]f;
	reg [15:0]g;
	reg [15:0]h;
	reg [2:0]sel;
	wire [15:0]out;
	
	mux_8way16bit_chip mux8way16bit(out, a, b, c, d, e, f, g, h, sel);

	initial begin
		$monitor("a: %b, b: %b, c: %b, d: %b, e: %b, f: %b, g: %b, h: %b, sel: %b,  out: %b", a, b, c, d, e, f, g, h, sel, out );	

		// initial conditions
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b000; #10

		// TEST case 1
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b000; #10
		// TEST case 2
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b001; #10
		// TEST case 3
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b010; #10
		// TEST case 4
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b011; #10
		// TEST case 5
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b100; #10
		// TEST case 6
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b101; #10
		// TEST case 7
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b110; #10
		// TEST case 8
		a = 16'b1000000000000000; b = 16'b0100000000000000; c = 16'b0010000000000000; d = 16'b0001000000000000;	e = 16'b0000100000000000; f = 16'b0000010000000000; g = 16'b0000001000000000; h = 16'b0000000100000000; sel = 3'b011; #10
		$finish;
	end

endmodule


