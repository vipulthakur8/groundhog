// One bit register

module bit(in load);
	input in, load;
endmodule
