module alu();
endmodule
